***** Spice Netlist for Cell 'Lab1' *****

************** Module Lab1 **************
v0 n0 gnd sin('0v' '4v' '1k') 
r0 n0 va 50 noisy=0 
r1 va vb 160k noisy=0 
c0 gnd vb 1.2f 


.end

